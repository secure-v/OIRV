//-----------------------interface signal---------------------------//
module BLACK_CELL(input Gi_k,
				  input Pi_k,
				  input Gk_1_j,
				  input Pk_1_j,
				  output Gi_j,
				  output Pi_j);
//////////////////////////////////////////////////////////////////////

//-----------------------internal signal----------------------------//
				  wire m;
//////////////////////////////////////////////////////////////////////

//-----------------------architecture-------------------------------//
				  and (Pi_j,Pi_k,Pk_1_j);

				  and (m,Pi_k,Gk_1_j);
				  or  (Gi_j,m,Gi_k);
//////////////////////////////////////////////////////////////////////
endmodule

