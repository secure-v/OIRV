module srt4_qds_table (
	input [6:0]        partial_sum,
	input [2:0]        d          ,
	output reg[2:0]    q          
);

	wire[9:0] index;
	assign index = {partial_sum, d};

	always@(*) begin
		case (index)
			10'd0: q = 3'b000;
			10'd1: q = 3'b000;
			10'd2: q = 3'b000;
			10'd3: q = 3'b000;
			10'd4: q = 3'b000;
			10'd5: q = 3'b000;
			10'd6: q = 3'b000;
			10'd7: q = 3'b000;
			10'd8: q = 3'b000;
			10'd9: q = 3'b000;
			10'd10: q = 3'b000;
			10'd11: q = 3'b000;
			10'd12: q = 3'b000;
			10'd13: q = 3'b000;
			10'd14: q = 3'b000;
			10'd15: q = 3'b000;
			10'd16: q = 3'b000;
			10'd17: q = 3'b000;
			10'd18: q = 3'b000;
			10'd19: q = 3'b000;
			10'd20: q = 3'b000;
			10'd21: q = 3'b000;
			10'd22: q = 3'b000;
			10'd23: q = 3'b000;
			10'd24: q = 3'b000;
			10'd25: q = 3'b000;
			10'd26: q = 3'b000;
			10'd27: q = 3'b000;
			10'd28: q = 3'b000;
			10'd29: q = 3'b000;
			10'd30: q = 3'b000;
			10'd31: q = 3'b000;
			10'd32: q = 3'b001;
			10'd33: q = 3'b001;
			10'd34: q = 3'b001;
			10'd35: q = 3'b001;
			10'd36: q = 3'b000;
			10'd37: q = 3'b000;
			10'd38: q = 3'b000;
			10'd39: q = 3'b000;
			10'd40: q = 3'b001;
			10'd41: q = 3'b001;
			10'd42: q = 3'b001;
			10'd43: q = 3'b001;
			10'd44: q = 3'b000;
			10'd45: q = 3'b000;
			10'd46: q = 3'b000;
			10'd47: q = 3'b000;
			10'd48: q = 3'b001;
			10'd49: q = 3'b001;
			10'd50: q = 3'b001;
			10'd51: q = 3'b001;
			10'd52: q = 3'b000;
			10'd53: q = 3'b000;
			10'd54: q = 3'b000;
			10'd55: q = 3'b000;
			10'd56: q = 3'b001;
			10'd57: q = 3'b001;
			10'd58: q = 3'b001;
			10'd59: q = 3'b001;
			10'd60: q = 3'b001;
			10'd61: q = 3'b001;
			10'd62: q = 3'b001;
			10'd63: q = 3'b001;
			10'd64: q = 3'b001;
			10'd65: q = 3'b001;
			10'd66: q = 3'b001;
			10'd67: q = 3'b001;
			10'd68: q = 3'b001;
			10'd69: q = 3'b001;
			10'd70: q = 3'b001;
			10'd71: q = 3'b001;
			10'd72: q = 3'b001;
			10'd73: q = 3'b001;
			10'd74: q = 3'b001;
			10'd75: q = 3'b001;
			10'd76: q = 3'b001;
			10'd77: q = 3'b001;
			10'd78: q = 3'b001;
			10'd79: q = 3'b001;
			10'd80: q = 3'b001;
			10'd81: q = 3'b001;
			10'd82: q = 3'b001;
			10'd83: q = 3'b001;
			10'd84: q = 3'b001;
			10'd85: q = 3'b001;
			10'd86: q = 3'b001;
			10'd87: q = 3'b001;
			10'd88: q = 3'b001;
			10'd89: q = 3'b001;
			10'd90: q = 3'b001;
			10'd91: q = 3'b001;
			10'd92: q = 3'b001;
			10'd93: q = 3'b001;
			10'd94: q = 3'b001;
			10'd95: q = 3'b001;
			10'd96: q = 3'b010;
			10'd97: q = 3'b001;
			10'd98: q = 3'b001;
			10'd99: q = 3'b001;
			10'd100: q = 3'b001;
			10'd101: q = 3'b001;
			10'd102: q = 3'b001;
			10'd103: q = 3'b001;
			10'd104: q = 3'b010;
			10'd105: q = 3'b001;
			10'd106: q = 3'b001;
			10'd107: q = 3'b001;
			10'd108: q = 3'b001;
			10'd109: q = 3'b001;
			10'd110: q = 3'b001;
			10'd111: q = 3'b001;
			10'd112: q = 3'b010;
			10'd113: q = 3'b010;
			10'd114: q = 3'b001;
			10'd115: q = 3'b001;
			10'd116: q = 3'b001;
			10'd117: q = 3'b001;
			10'd118: q = 3'b001;
			10'd119: q = 3'b001;
			10'd120: q = 3'b010;
			10'd121: q = 3'b010;
			10'd122: q = 3'b010;
			10'd123: q = 3'b001;
			10'd124: q = 3'b001;
			10'd125: q = 3'b001;
			10'd126: q = 3'b001;
			10'd127: q = 3'b001;
			10'd128: q = 3'b010;
			10'd129: q = 3'b010;
			10'd130: q = 3'b010;
			10'd131: q = 3'b001;
			10'd132: q = 3'b001;
			10'd133: q = 3'b001;
			10'd134: q = 3'b001;
			10'd135: q = 3'b001;
			10'd136: q = 3'b010;
			10'd137: q = 3'b010;
			10'd138: q = 3'b010;
			10'd139: q = 3'b010;
			10'd140: q = 3'b001;
			10'd141: q = 3'b001;
			10'd142: q = 3'b001;
			10'd143: q = 3'b001;
			10'd144: q = 3'b010;
			10'd145: q = 3'b010;
			10'd146: q = 3'b010;
			10'd147: q = 3'b010;
			10'd148: q = 3'b001;
			10'd149: q = 3'b001;
			10'd150: q = 3'b001;
			10'd151: q = 3'b001;
			10'd152: q = 3'b010;
			10'd153: q = 3'b010;
			10'd154: q = 3'b010;
			10'd155: q = 3'b010;
			10'd156: q = 3'b010;
			10'd157: q = 3'b010;
			10'd158: q = 3'b001;
			10'd159: q = 3'b001;
			10'd160: q = 3'b010;
			10'd161: q = 3'b010;
			10'd162: q = 3'b010;
			10'd163: q = 3'b010;
			10'd164: q = 3'b010;
			10'd165: q = 3'b010;
			10'd166: q = 3'b001;
			10'd167: q = 3'b001;
			10'd168: q = 3'b010;
			10'd169: q = 3'b010;
			10'd170: q = 3'b010;
			10'd171: q = 3'b010;
			10'd172: q = 3'b010;
			10'd173: q = 3'b010;
			10'd174: q = 3'b010;
			10'd175: q = 3'b001;
			10'd176: q = 3'b010;
			10'd177: q = 3'b010;
			10'd178: q = 3'b010;
			10'd179: q = 3'b010;
			10'd180: q = 3'b010;
			10'd181: q = 3'b010;
			10'd182: q = 3'b010;
			10'd183: q = 3'b001;
			10'd184: q = 3'b010;
			10'd185: q = 3'b010;
			10'd186: q = 3'b010;
			10'd187: q = 3'b010;
			10'd188: q = 3'b010;
			10'd189: q = 3'b010;
			10'd190: q = 3'b010;
			10'd191: q = 3'b010;
			10'd192: q = 3'b010;
			10'd193: q = 3'b010;
			10'd194: q = 3'b010;
			10'd195: q = 3'b010;
			10'd196: q = 3'b010;
			10'd197: q = 3'b010;
			10'd198: q = 3'b010;
			10'd199: q = 3'b010;
			10'd200: q = 3'b010;
			10'd201: q = 3'b010;
			10'd202: q = 3'b010;
			10'd203: q = 3'b010;
			10'd204: q = 3'b010;
			10'd205: q = 3'b010;
			10'd206: q = 3'b010;
			10'd207: q = 3'b010;
			10'd208: q = 3'b010;
			10'd209: q = 3'b010;
			10'd210: q = 3'b010;
			10'd211: q = 3'b010;
			10'd212: q = 3'b010;
			10'd213: q = 3'b010;
			10'd214: q = 3'b010;
			10'd215: q = 3'b010;
			10'd216: q = 3'b010;
			10'd217: q = 3'b010;
			10'd218: q = 3'b010;
			10'd219: q = 3'b010;
			10'd220: q = 3'b010;
			10'd221: q = 3'b010;
			10'd222: q = 3'b010;
			10'd223: q = 3'b010;
			10'd224: q = 3'b010;
			10'd225: q = 3'b010;
			10'd226: q = 3'b010;
			10'd227: q = 3'b010;
			10'd228: q = 3'b010;
			10'd229: q = 3'b010;
			10'd230: q = 3'b010;
			10'd231: q = 3'b010;
			10'd232: q = 3'b010;
			10'd233: q = 3'b010;
			10'd234: q = 3'b010;
			10'd235: q = 3'b010;
			10'd236: q = 3'b010;
			10'd237: q = 3'b010;
			10'd238: q = 3'b010;
			10'd239: q = 3'b010;
			10'd240: q = 3'b010;
			10'd241: q = 3'b010;
			10'd242: q = 3'b010;
			10'd243: q = 3'b010;
			10'd244: q = 3'b010;
			10'd245: q = 3'b010;
			10'd246: q = 3'b010;
			10'd247: q = 3'b010;
			10'd248: q = 3'b010;
			10'd249: q = 3'b010;
			10'd250: q = 3'b010;
			10'd251: q = 3'b010;
			10'd252: q = 3'b010;
			10'd253: q = 3'b010;
			10'd254: q = 3'b010;
			10'd255: q = 3'b010;
			10'd256: q = 3'b010;
			10'd257: q = 3'b010;
			10'd258: q = 3'b010;
			10'd259: q = 3'b010;
			10'd260: q = 3'b010;
			10'd261: q = 3'b010;
			10'd262: q = 3'b010;
			10'd263: q = 3'b010;
			10'd264: q = 3'b010;
			10'd265: q = 3'b010;
			10'd266: q = 3'b010;
			10'd267: q = 3'b010;
			10'd268: q = 3'b010;
			10'd269: q = 3'b010;
			10'd270: q = 3'b010;
			10'd271: q = 3'b010;
			10'd272: q = 3'b010;
			10'd273: q = 3'b010;
			10'd274: q = 3'b010;
			10'd275: q = 3'b010;
			10'd276: q = 3'b010;
			10'd277: q = 3'b010;
			10'd278: q = 3'b010;
			10'd279: q = 3'b010;
			10'd280: q = 3'b010;
			10'd281: q = 3'b010;
			10'd282: q = 3'b010;
			10'd283: q = 3'b010;
			10'd284: q = 3'b010;
			10'd285: q = 3'b010;
			10'd286: q = 3'b010;
			10'd287: q = 3'b010;
			10'd288: q = 3'b010;
			10'd289: q = 3'b010;
			10'd290: q = 3'b010;
			10'd291: q = 3'b010;
			10'd292: q = 3'b010;
			10'd293: q = 3'b010;
			10'd294: q = 3'b010;
			10'd295: q = 3'b010;
			10'd296: q = 3'b010;
			10'd297: q = 3'b010;
			10'd298: q = 3'b010;
			10'd299: q = 3'b010;
			10'd300: q = 3'b010;
			10'd301: q = 3'b010;
			10'd302: q = 3'b010;
			10'd303: q = 3'b010;
			10'd304: q = 3'b010;
			10'd305: q = 3'b010;
			10'd306: q = 3'b010;
			10'd307: q = 3'b010;
			10'd308: q = 3'b010;
			10'd309: q = 3'b010;
			10'd310: q = 3'b010;
			10'd311: q = 3'b010;
			10'd312: q = 3'b010;
			10'd313: q = 3'b010;
			10'd314: q = 3'b010;
			10'd315: q = 3'b010;
			10'd316: q = 3'b010;
			10'd317: q = 3'b010;
			10'd318: q = 3'b010;
			10'd319: q = 3'b010;
			10'd320: q = 3'b010;
			10'd321: q = 3'b010;
			10'd322: q = 3'b010;
			10'd323: q = 3'b010;
			10'd324: q = 3'b010;
			10'd325: q = 3'b010;
			10'd326: q = 3'b010;
			10'd327: q = 3'b010;
			10'd328: q = 3'b010;
			10'd329: q = 3'b010;
			10'd330: q = 3'b010;
			10'd331: q = 3'b010;
			10'd332: q = 3'b010;
			10'd333: q = 3'b010;
			10'd334: q = 3'b010;
			10'd335: q = 3'b010;
			10'd336: q = 3'b010;
			10'd337: q = 3'b010;
			10'd338: q = 3'b010;
			10'd339: q = 3'b010;
			10'd340: q = 3'b010;
			10'd341: q = 3'b010;
			10'd342: q = 3'b010;
			10'd343: q = 3'b010;
			10'd344: q = 3'b010;
			10'd345: q = 3'b010;
			10'd346: q = 3'b010;
			10'd347: q = 3'b010;
			10'd348: q = 3'b010;
			10'd349: q = 3'b010;
			10'd350: q = 3'b010;
			10'd351: q = 3'b010;
			10'd352: q = 3'b010;
			10'd353: q = 3'b010;
			10'd354: q = 3'b010;
			10'd355: q = 3'b010;
			10'd356: q = 3'b010;
			10'd357: q = 3'b010;
			10'd358: q = 3'b010;
			10'd359: q = 3'b010;
			10'd360: q = 3'b010;
			10'd361: q = 3'b010;
			10'd362: q = 3'b010;
			10'd363: q = 3'b010;
			10'd364: q = 3'b010;
			10'd365: q = 3'b010;
			10'd366: q = 3'b010;
			10'd367: q = 3'b010;
			10'd368: q = 3'b010;
			10'd369: q = 3'b010;
			10'd370: q = 3'b010;
			10'd371: q = 3'b010;
			10'd372: q = 3'b010;
			10'd373: q = 3'b010;
			10'd374: q = 3'b010;
			10'd375: q = 3'b010;
			10'd376: q = 3'b010;
			10'd377: q = 3'b010;
			10'd378: q = 3'b010;
			10'd379: q = 3'b010;
			10'd380: q = 3'b010;
			10'd381: q = 3'b010;
			10'd382: q = 3'b010;
			10'd383: q = 3'b010;
			10'd384: q = 3'b010;
			10'd385: q = 3'b010;
			10'd386: q = 3'b010;
			10'd387: q = 3'b010;
			10'd388: q = 3'b010;
			10'd389: q = 3'b010;
			10'd390: q = 3'b010;
			10'd391: q = 3'b010;
			10'd392: q = 3'b010;
			10'd393: q = 3'b010;
			10'd394: q = 3'b010;
			10'd395: q = 3'b010;
			10'd396: q = 3'b010;
			10'd397: q = 3'b010;
			10'd398: q = 3'b010;
			10'd399: q = 3'b010;
			10'd400: q = 3'b010;
			10'd401: q = 3'b010;
			10'd402: q = 3'b010;
			10'd403: q = 3'b010;
			10'd404: q = 3'b010;
			10'd405: q = 3'b010;
			10'd406: q = 3'b010;
			10'd407: q = 3'b010;
			10'd408: q = 3'b010;
			10'd409: q = 3'b010;
			10'd410: q = 3'b010;
			10'd411: q = 3'b010;
			10'd412: q = 3'b010;
			10'd413: q = 3'b010;
			10'd414: q = 3'b010;
			10'd415: q = 3'b010;
			10'd416: q = 3'b010;
			10'd417: q = 3'b010;
			10'd418: q = 3'b010;
			10'd419: q = 3'b010;
			10'd420: q = 3'b010;
			10'd421: q = 3'b010;
			10'd422: q = 3'b010;
			10'd423: q = 3'b010;
			10'd424: q = 3'b010;
			10'd425: q = 3'b010;
			10'd426: q = 3'b010;
			10'd427: q = 3'b010;
			10'd428: q = 3'b010;
			10'd429: q = 3'b010;
			10'd430: q = 3'b010;
			10'd431: q = 3'b010;
			10'd432: q = 3'b010;
			10'd433: q = 3'b010;
			10'd434: q = 3'b010;
			10'd435: q = 3'b010;
			10'd436: q = 3'b010;
			10'd437: q = 3'b010;
			10'd438: q = 3'b010;
			10'd439: q = 3'b010;
			10'd440: q = 3'b010;
			10'd441: q = 3'b010;
			10'd442: q = 3'b010;
			10'd443: q = 3'b010;
			10'd444: q = 3'b010;
			10'd445: q = 3'b010;
			10'd446: q = 3'b010;
			10'd447: q = 3'b010;
			10'd448: q = 3'b010;
			10'd449: q = 3'b010;
			10'd450: q = 3'b010;
			10'd451: q = 3'b010;
			10'd452: q = 3'b010;
			10'd453: q = 3'b010;
			10'd454: q = 3'b010;
			10'd455: q = 3'b010;
			10'd456: q = 3'b010;
			10'd457: q = 3'b010;
			10'd458: q = 3'b010;
			10'd459: q = 3'b010;
			10'd460: q = 3'b010;
			10'd461: q = 3'b010;
			10'd462: q = 3'b010;
			10'd463: q = 3'b010;
			10'd464: q = 3'b010;
			10'd465: q = 3'b010;
			10'd466: q = 3'b010;
			10'd467: q = 3'b010;
			10'd468: q = 3'b010;
			10'd469: q = 3'b010;
			10'd470: q = 3'b010;
			10'd471: q = 3'b010;
			10'd472: q = 3'b010;
			10'd473: q = 3'b010;
			10'd474: q = 3'b010;
			10'd475: q = 3'b010;
			10'd476: q = 3'b010;
			10'd477: q = 3'b010;
			10'd478: q = 3'b010;
			10'd479: q = 3'b010;
			10'd480: q = 3'b010;
			10'd481: q = 3'b010;
			10'd482: q = 3'b010;
			10'd483: q = 3'b010;
			10'd484: q = 3'b010;
			10'd485: q = 3'b010;
			10'd486: q = 3'b010;
			10'd487: q = 3'b010;
			10'd488: q = 3'b010;
			10'd489: q = 3'b010;
			10'd490: q = 3'b010;
			10'd491: q = 3'b010;
			10'd492: q = 3'b010;
			10'd493: q = 3'b010;
			10'd494: q = 3'b010;
			10'd495: q = 3'b010;
			10'd496: q = 3'b010;
			10'd497: q = 3'b010;
			10'd498: q = 3'b010;
			10'd499: q = 3'b010;
			10'd500: q = 3'b010;
			10'd501: q = 3'b010;
			10'd502: q = 3'b010;
			10'd503: q = 3'b010;
			10'd504: q = 3'b010;
			10'd505: q = 3'b010;
			10'd506: q = 3'b010;
			10'd507: q = 3'b010;
			10'd508: q = 3'b010;
			10'd509: q = 3'b010;
			10'd510: q = 3'b010;
			10'd511: q = 3'b010;
			10'd512: q = 3'b110;
			10'd513: q = 3'b110;
			10'd514: q = 3'b110;
			10'd515: q = 3'b110;
			10'd516: q = 3'b110;
			10'd517: q = 3'b110;
			10'd518: q = 3'b110;
			10'd519: q = 3'b110;
			10'd520: q = 3'b110;
			10'd521: q = 3'b110;
			10'd522: q = 3'b110;
			10'd523: q = 3'b110;
			10'd524: q = 3'b110;
			10'd525: q = 3'b110;
			10'd526: q = 3'b110;
			10'd527: q = 3'b110;
			10'd528: q = 3'b110;
			10'd529: q = 3'b110;
			10'd530: q = 3'b110;
			10'd531: q = 3'b110;
			10'd532: q = 3'b110;
			10'd533: q = 3'b110;
			10'd534: q = 3'b110;
			10'd535: q = 3'b110;
			10'd536: q = 3'b110;
			10'd537: q = 3'b110;
			10'd538: q = 3'b110;
			10'd539: q = 3'b110;
			10'd540: q = 3'b110;
			10'd541: q = 3'b110;
			10'd542: q = 3'b110;
			10'd543: q = 3'b110;
			10'd544: q = 3'b110;
			10'd545: q = 3'b110;
			10'd546: q = 3'b110;
			10'd547: q = 3'b110;
			10'd548: q = 3'b110;
			10'd549: q = 3'b110;
			10'd550: q = 3'b110;
			10'd551: q = 3'b110;
			10'd552: q = 3'b110;
			10'd553: q = 3'b110;
			10'd554: q = 3'b110;
			10'd555: q = 3'b110;
			10'd556: q = 3'b110;
			10'd557: q = 3'b110;
			10'd558: q = 3'b110;
			10'd559: q = 3'b110;
			10'd560: q = 3'b110;
			10'd561: q = 3'b110;
			10'd562: q = 3'b110;
			10'd563: q = 3'b110;
			10'd564: q = 3'b110;
			10'd565: q = 3'b110;
			10'd566: q = 3'b110;
			10'd567: q = 3'b110;
			10'd568: q = 3'b110;
			10'd569: q = 3'b110;
			10'd570: q = 3'b110;
			10'd571: q = 3'b110;
			10'd572: q = 3'b110;
			10'd573: q = 3'b110;
			10'd574: q = 3'b110;
			10'd575: q = 3'b110;
			10'd576: q = 3'b110;
			10'd577: q = 3'b110;
			10'd578: q = 3'b110;
			10'd579: q = 3'b110;
			10'd580: q = 3'b110;
			10'd581: q = 3'b110;
			10'd582: q = 3'b110;
			10'd583: q = 3'b110;
			10'd584: q = 3'b110;
			10'd585: q = 3'b110;
			10'd586: q = 3'b110;
			10'd587: q = 3'b110;
			10'd588: q = 3'b110;
			10'd589: q = 3'b110;
			10'd590: q = 3'b110;
			10'd591: q = 3'b110;
			10'd592: q = 3'b110;
			10'd593: q = 3'b110;
			10'd594: q = 3'b110;
			10'd595: q = 3'b110;
			10'd596: q = 3'b110;
			10'd597: q = 3'b110;
			10'd598: q = 3'b110;
			10'd599: q = 3'b110;
			10'd600: q = 3'b110;
			10'd601: q = 3'b110;
			10'd602: q = 3'b110;
			10'd603: q = 3'b110;
			10'd604: q = 3'b110;
			10'd605: q = 3'b110;
			10'd606: q = 3'b110;
			10'd607: q = 3'b110;
			10'd608: q = 3'b110;
			10'd609: q = 3'b110;
			10'd610: q = 3'b110;
			10'd611: q = 3'b110;
			10'd612: q = 3'b110;
			10'd613: q = 3'b110;
			10'd614: q = 3'b110;
			10'd615: q = 3'b110;
			10'd616: q = 3'b110;
			10'd617: q = 3'b110;
			10'd618: q = 3'b110;
			10'd619: q = 3'b110;
			10'd620: q = 3'b110;
			10'd621: q = 3'b110;
			10'd622: q = 3'b110;
			10'd623: q = 3'b110;
			10'd624: q = 3'b110;
			10'd625: q = 3'b110;
			10'd626: q = 3'b110;
			10'd627: q = 3'b110;
			10'd628: q = 3'b110;
			10'd629: q = 3'b110;
			10'd630: q = 3'b110;
			10'd631: q = 3'b110;
			10'd632: q = 3'b110;
			10'd633: q = 3'b110;
			10'd634: q = 3'b110;
			10'd635: q = 3'b110;
			10'd636: q = 3'b110;
			10'd637: q = 3'b110;
			10'd638: q = 3'b110;
			10'd639: q = 3'b110;
			10'd640: q = 3'b110;
			10'd641: q = 3'b110;
			10'd642: q = 3'b110;
			10'd643: q = 3'b110;
			10'd644: q = 3'b110;
			10'd645: q = 3'b110;
			10'd646: q = 3'b110;
			10'd647: q = 3'b110;
			10'd648: q = 3'b110;
			10'd649: q = 3'b110;
			10'd650: q = 3'b110;
			10'd651: q = 3'b110;
			10'd652: q = 3'b110;
			10'd653: q = 3'b110;
			10'd654: q = 3'b110;
			10'd655: q = 3'b110;
			10'd656: q = 3'b110;
			10'd657: q = 3'b110;
			10'd658: q = 3'b110;
			10'd659: q = 3'b110;
			10'd660: q = 3'b110;
			10'd661: q = 3'b110;
			10'd662: q = 3'b110;
			10'd663: q = 3'b110;
			10'd664: q = 3'b110;
			10'd665: q = 3'b110;
			10'd666: q = 3'b110;
			10'd667: q = 3'b110;
			10'd668: q = 3'b110;
			10'd669: q = 3'b110;
			10'd670: q = 3'b110;
			10'd671: q = 3'b110;
			10'd672: q = 3'b110;
			10'd673: q = 3'b110;
			10'd674: q = 3'b110;
			10'd675: q = 3'b110;
			10'd676: q = 3'b110;
			10'd677: q = 3'b110;
			10'd678: q = 3'b110;
			10'd679: q = 3'b110;
			10'd680: q = 3'b110;
			10'd681: q = 3'b110;
			10'd682: q = 3'b110;
			10'd683: q = 3'b110;
			10'd684: q = 3'b110;
			10'd685: q = 3'b110;
			10'd686: q = 3'b110;
			10'd687: q = 3'b110;
			10'd688: q = 3'b110;
			10'd689: q = 3'b110;
			10'd690: q = 3'b110;
			10'd691: q = 3'b110;
			10'd692: q = 3'b110;
			10'd693: q = 3'b110;
			10'd694: q = 3'b110;
			10'd695: q = 3'b110;
			10'd696: q = 3'b110;
			10'd697: q = 3'b110;
			10'd698: q = 3'b110;
			10'd699: q = 3'b110;
			10'd700: q = 3'b110;
			10'd701: q = 3'b110;
			10'd702: q = 3'b110;
			10'd703: q = 3'b110;
			10'd704: q = 3'b110;
			10'd705: q = 3'b110;
			10'd706: q = 3'b110;
			10'd707: q = 3'b110;
			10'd708: q = 3'b110;
			10'd709: q = 3'b110;
			10'd710: q = 3'b110;
			10'd711: q = 3'b110;
			10'd712: q = 3'b110;
			10'd713: q = 3'b110;
			10'd714: q = 3'b110;
			10'd715: q = 3'b110;
			10'd716: q = 3'b110;
			10'd717: q = 3'b110;
			10'd718: q = 3'b110;
			10'd719: q = 3'b110;
			10'd720: q = 3'b110;
			10'd721: q = 3'b110;
			10'd722: q = 3'b110;
			10'd723: q = 3'b110;
			10'd724: q = 3'b110;
			10'd725: q = 3'b110;
			10'd726: q = 3'b110;
			10'd727: q = 3'b110;
			10'd728: q = 3'b110;
			10'd729: q = 3'b110;
			10'd730: q = 3'b110;
			10'd731: q = 3'b110;
			10'd732: q = 3'b110;
			10'd733: q = 3'b110;
			10'd734: q = 3'b110;
			10'd735: q = 3'b110;
			10'd736: q = 3'b110;
			10'd737: q = 3'b110;
			10'd738: q = 3'b110;
			10'd739: q = 3'b110;
			10'd740: q = 3'b110;
			10'd741: q = 3'b110;
			10'd742: q = 3'b110;
			10'd743: q = 3'b110;
			10'd744: q = 3'b110;
			10'd745: q = 3'b110;
			10'd746: q = 3'b110;
			10'd747: q = 3'b110;
			10'd748: q = 3'b110;
			10'd749: q = 3'b110;
			10'd750: q = 3'b110;
			10'd751: q = 3'b110;
			10'd752: q = 3'b110;
			10'd753: q = 3'b110;
			10'd754: q = 3'b110;
			10'd755: q = 3'b110;
			10'd756: q = 3'b110;
			10'd757: q = 3'b110;
			10'd758: q = 3'b110;
			10'd759: q = 3'b110;
			10'd760: q = 3'b110;
			10'd761: q = 3'b110;
			10'd762: q = 3'b110;
			10'd763: q = 3'b110;
			10'd764: q = 3'b110;
			10'd765: q = 3'b110;
			10'd766: q = 3'b110;
			10'd767: q = 3'b110;
			10'd768: q = 3'b110;
			10'd769: q = 3'b110;
			10'd770: q = 3'b110;
			10'd771: q = 3'b110;
			10'd772: q = 3'b110;
			10'd773: q = 3'b110;
			10'd774: q = 3'b110;
			10'd775: q = 3'b110;
			10'd776: q = 3'b110;
			10'd777: q = 3'b110;
			10'd778: q = 3'b110;
			10'd779: q = 3'b110;
			10'd780: q = 3'b110;
			10'd781: q = 3'b110;
			10'd782: q = 3'b110;
			10'd783: q = 3'b110;
			10'd784: q = 3'b110;
			10'd785: q = 3'b110;
			10'd786: q = 3'b110;
			10'd787: q = 3'b110;
			10'd788: q = 3'b110;
			10'd789: q = 3'b110;
			10'd790: q = 3'b110;
			10'd791: q = 3'b110;
			10'd792: q = 3'b110;
			10'd793: q = 3'b110;
			10'd794: q = 3'b110;
			10'd795: q = 3'b110;
			10'd796: q = 3'b110;
			10'd797: q = 3'b110;
			10'd798: q = 3'b110;
			10'd799: q = 3'b110;
			10'd800: q = 3'b110;
			10'd801: q = 3'b110;
			10'd802: q = 3'b110;
			10'd803: q = 3'b110;
			10'd804: q = 3'b110;
			10'd805: q = 3'b110;
			10'd806: q = 3'b110;
			10'd807: q = 3'b110;
			10'd808: q = 3'b110;
			10'd809: q = 3'b110;
			10'd810: q = 3'b110;
			10'd811: q = 3'b110;
			10'd812: q = 3'b110;
			10'd813: q = 3'b110;
			10'd814: q = 3'b110;
			10'd815: q = 3'b110;
			10'd816: q = 3'b110;
			10'd817: q = 3'b110;
			10'd818: q = 3'b110;
			10'd819: q = 3'b110;
			10'd820: q = 3'b110;
			10'd821: q = 3'b110;
			10'd822: q = 3'b110;
			10'd823: q = 3'b110;
			10'd824: q = 3'b110;
			10'd825: q = 3'b110;
			10'd826: q = 3'b110;
			10'd827: q = 3'b110;
			10'd828: q = 3'b110;
			10'd829: q = 3'b110;
			10'd830: q = 3'b110;
			10'd831: q = 3'b110;
			10'd832: q = 3'b110;
			10'd833: q = 3'b110;
			10'd834: q = 3'b110;
			10'd835: q = 3'b110;
			10'd836: q = 3'b110;
			10'd837: q = 3'b110;
			10'd838: q = 3'b110;
			10'd839: q = 3'b110;
			10'd840: q = 3'b110;
			10'd841: q = 3'b110;
			10'd842: q = 3'b110;
			10'd843: q = 3'b110;
			10'd844: q = 3'b110;
			10'd845: q = 3'b110;
			10'd846: q = 3'b110;
			10'd847: q = 3'b110;
			10'd848: q = 3'b110;
			10'd849: q = 3'b110;
			10'd850: q = 3'b110;
			10'd851: q = 3'b110;
			10'd852: q = 3'b110;
			10'd853: q = 3'b110;
			10'd854: q = 3'b101;
			10'd855: q = 3'b101;
			10'd856: q = 3'b110;
			10'd857: q = 3'b110;
			10'd858: q = 3'b110;
			10'd859: q = 3'b110;
			10'd860: q = 3'b110;
			10'd861: q = 3'b110;
			10'd862: q = 3'b101;
			10'd863: q = 3'b101;
			10'd864: q = 3'b110;
			10'd865: q = 3'b110;
			10'd866: q = 3'b110;
			10'd867: q = 3'b110;
			10'd868: q = 3'b101;
			10'd869: q = 3'b101;
			10'd870: q = 3'b101;
			10'd871: q = 3'b101;
			10'd872: q = 3'b110;
			10'd873: q = 3'b110;
			10'd874: q = 3'b110;
			10'd875: q = 3'b110;
			10'd876: q = 3'b101;
			10'd877: q = 3'b101;
			10'd878: q = 3'b101;
			10'd879: q = 3'b101;
			10'd880: q = 3'b110;
			10'd881: q = 3'b110;
			10'd882: q = 3'b110;
			10'd883: q = 3'b101;
			10'd884: q = 3'b101;
			10'd885: q = 3'b101;
			10'd886: q = 3'b101;
			10'd887: q = 3'b101;
			10'd888: q = 3'b110;
			10'd889: q = 3'b110;
			10'd890: q = 3'b110;
			10'd891: q = 3'b101;
			10'd892: q = 3'b101;
			10'd893: q = 3'b101;
			10'd894: q = 3'b101;
			10'd895: q = 3'b101;
			10'd896: q = 3'b110;
			10'd897: q = 3'b110;
			10'd898: q = 3'b101;
			10'd899: q = 3'b101;
			10'd900: q = 3'b101;
			10'd901: q = 3'b101;
			10'd902: q = 3'b101;
			10'd903: q = 3'b101;
			10'd904: q = 3'b110;
			10'd905: q = 3'b110;
			10'd906: q = 3'b101;
			10'd907: q = 3'b101;
			10'd908: q = 3'b101;
			10'd909: q = 3'b101;
			10'd910: q = 3'b101;
			10'd911: q = 3'b101;
			10'd912: q = 3'b110;
			10'd913: q = 3'b101;
			10'd914: q = 3'b101;
			10'd915: q = 3'b101;
			10'd916: q = 3'b101;
			10'd917: q = 3'b101;
			10'd918: q = 3'b101;
			10'd919: q = 3'b101;
			10'd920: q = 3'b101;
			10'd921: q = 3'b101;
			10'd922: q = 3'b101;
			10'd923: q = 3'b101;
			10'd924: q = 3'b101;
			10'd925: q = 3'b101;
			10'd926: q = 3'b101;
			10'd927: q = 3'b101;
			10'd928: q = 3'b101;
			10'd929: q = 3'b101;
			10'd930: q = 3'b101;
			10'd931: q = 3'b101;
			10'd932: q = 3'b101;
			10'd933: q = 3'b101;
			10'd934: q = 3'b101;
			10'd935: q = 3'b101;
			10'd936: q = 3'b101;
			10'd937: q = 3'b101;
			10'd938: q = 3'b101;
			10'd939: q = 3'b101;
			10'd940: q = 3'b101;
			10'd941: q = 3'b101;
			10'd942: q = 3'b101;
			10'd943: q = 3'b101;
			10'd944: q = 3'b101;
			10'd945: q = 3'b101;
			10'd946: q = 3'b101;
			10'd947: q = 3'b101;
			10'd948: q = 3'b101;
			10'd949: q = 3'b101;
			10'd950: q = 3'b101;
			10'd951: q = 3'b101;
			10'd952: q = 3'b101;
			10'd953: q = 3'b101;
			10'd954: q = 3'b101;
			10'd955: q = 3'b101;
			10'd956: q = 3'b101;
			10'd957: q = 3'b101;
			10'd958: q = 3'b101;
			10'd959: q = 3'b101;
			10'd960: q = 3'b101;
			10'd961: q = 3'b101;
			10'd962: q = 3'b101;
			10'd963: q = 3'b101;
			10'd964: q = 3'b101;
			10'd965: q = 3'b101;
			10'd966: q = 3'b101;
			10'd967: q = 3'b101;
			10'd968: q = 3'b101;
			10'd969: q = 3'b101;
			10'd970: q = 3'b101;
			10'd971: q = 3'b101;
			10'd972: q = 3'b101;
			10'd973: q = 3'b101;
			10'd974: q = 3'b101;
			10'd975: q = 3'b101;
			10'd976: q = 3'b101;
			10'd977: q = 3'b101;
			10'd978: q = 3'b101;
			10'd979: q = 3'b101;
			10'd980: q = 3'b000;
			10'd981: q = 3'b000;
			10'd982: q = 3'b000;
			10'd983: q = 3'b000;
			10'd984: q = 3'b000;
			10'd985: q = 3'b000;
			10'd986: q = 3'b000;
			10'd987: q = 3'b000;
			10'd988: q = 3'b000;
			10'd989: q = 3'b000;
			10'd990: q = 3'b000;
			10'd991: q = 3'b000;
			10'd992: q = 3'b000;
			10'd993: q = 3'b000;
			10'd994: q = 3'b000;
			10'd995: q = 3'b000;
			10'd996: q = 3'b000;
			10'd997: q = 3'b000;
			10'd998: q = 3'b000;
			10'd999: q = 3'b000;
			10'd1000: q = 3'b000;
			10'd1001: q = 3'b000;
			10'd1002: q = 3'b000;
			10'd1003: q = 3'b000;
			10'd1004: q = 3'b000;
			10'd1005: q = 3'b000;
			10'd1006: q = 3'b000;
			10'd1007: q = 3'b000;
			10'd1008: q = 3'b000;
			10'd1009: q = 3'b000;
			10'd1010: q = 3'b000;
			10'd1011: q = 3'b000;
			10'd1012: q = 3'b000;
			10'd1013: q = 3'b000;
			10'd1014: q = 3'b000;
			10'd1015: q = 3'b000;
			10'd1016: q = 3'b000;
			10'd1017: q = 3'b000;
			10'd1018: q = 3'b000;
			10'd1019: q = 3'b000;
			10'd1020: q = 3'b000;
			10'd1021: q = 3'b000;
			10'd1022: q = 3'b000;
			10'd1023: q = 3'b000;
			default: q = 3'b000;
		endcase
	end

endmodule