//-----------------------interface signal---------------------------//
module GRAY_CELL(input Gi_k,
				 input Pi_k,
				 input Gk_1_j,
				 output Gi_j);
//////////////////////////////////////////////////////////////////////

//-----------------------internal signal----------------------------//
				 wire m;
//////////////////////////////////////////////////////////////////////

//-----------------------architecture-------------------------------//
				 and (m,Pi_k,Gk_1_j);
				 or  (Gi_j,m,Gi_k);
//////////////////////////////////////////////////////////////////////
endmodule

